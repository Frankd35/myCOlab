module branch_solver (
    ports
);
    
endmodule