`timescale 1ns / 1ps

module ClkDiv();

endmodule